magic
tech sky130A
timestamp 1609431327
<< end >>
