magic
tech sky130A
timestamp 1609332184
<< error_p >>
rect -38 -30 0 25
rect 15 -30 55 25
<< nmos >>
rect 0 -30 15 25
<< ndiff >>
rect -38 15 0 25
rect -38 -20 -33 15
rect -10 -20 0 15
rect -38 -30 0 -20
rect 15 15 55 25
rect 15 -20 30 15
rect 50 -20 55 15
rect 15 -30 55 -20
<< ndiffc >>
rect -33 -20 -10 15
rect 30 -20 50 15
<< poly >>
rect -25 70 15 80
rect -25 50 -20 70
rect 0 50 15 70
rect -25 40 15 50
rect 69 72 108 88
rect 640 87 679 91
rect 69 53 81 72
rect 100 53 108 72
rect 69 41 108 53
rect 634 81 679 87
rect 634 49 643 81
rect 667 49 679 81
rect 634 42 679 49
rect 634 41 672 42
rect -20 35 15 40
rect 0 25 15 35
rect 0 -45 15 -30
<< polycont >>
rect -20 50 0 70
rect 81 53 100 72
rect 643 49 667 81
<< npolyres >>
rect 108 41 634 87
<< locali >>
rect 30 87 70 89
rect -45 70 10 75
rect -45 50 -20 70
rect 0 50 10 70
rect -45 45 10 50
rect 30 72 100 87
rect 639 81 682 91
rect 30 53 81 72
rect 100 53 102 72
rect 30 41 100 53
rect 639 49 643 81
rect 667 49 682 81
rect -33 15 -10 25
rect -33 -65 -10 -20
rect 30 15 70 41
rect 639 37 682 49
rect 50 -20 70 15
rect 30 -33 70 -20
<< viali >>
rect -33 -87 -10 -65
<< metal1 >>
rect -59 -65 5 -41
rect -59 -87 -33 -65
rect -10 -87 5 -65
rect -59 -110 5 -87
<< labels >>
rlabel locali -45 45 -25 75 1 gate
rlabel metal1 -55 -105 -36 -71 1 VGND
rlabel ndiffc 30 -20 50 15 1 out
rlabel polycont 643 49 667 81 1 VPWR
<< end >>
