MOSFET Simulation
* this file edited to remove everything not in tt lib
.lib "./sky130_fd_pr/models/sky130.lib.spice" tt

* instantiate the inverter
Xmosfet VPWR A Y VGND VGND X0

.subckt X0 VPWR gate out VGND VSUBS
* NGSPICE file created from mosfet.ext - technology: sky130A


* Top level circuit mosfet

X0 out gate VGND VSUBS sky130_fd_pr__nfet_01v8 w=550000u l=150000u
R0 out VPWR sky130_fd_pr__res_generic_po w=460000u l=5.26e+06u
C0 out gate 0.07fF
C1 out VGND 0.05fF
C2 VGND gate 0.04fF
C3 VGND VSUBS 0.19fF
C4 VPWR VSUBS 0.19fF
C5 out VSUBS 0.11fF
C6 gate VSUBS 0.18fF


.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
Vin A VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10e-12 2e-09 0e-00

.control
run
set color0 = white
set color1 = black
plot A Y
plot i(Vdd)
.endc

.end
