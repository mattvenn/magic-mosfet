magic
tech sky130A
timestamp 1609431286
<< nmos >>
rect 40 0 55 65
<< ndiff >>
rect 0 0 40 65
rect 55 0 95 65
<< poly >>
rect 40 65 55 105
rect 40 -45 55 0
<< labels >>
rlabel ndiff 72 19 86 52 1 drain
rlabel ndiff 6 17 20 50 1 source
rlabel poly 40 -45 55 -10 1 gate
<< end >>
