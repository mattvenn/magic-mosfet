MOSFET Simulation
* this file edited to remove everything not in tt lib
.lib "./sky130_fd_pr/models/sky130.lib.spice" tt
.inc "sky130_fd_pr__res_generic_po.spice"

* instantiate the inverter
Xmosfet DRAIN GATE VGND VGND X0

.subckt X0 drain gate source VSUBS
* NGSPICE file created from mosfet.ext - technology: sky130A


* Top level circuit mosfet

X0 drain gate source VSUBS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
C0 drain source 0.06fF
C1 gate source 0.20fF
C2 drain VSUBS 0.15fF
C3 source VSUBS 0.15fF
C4 gate VSUBS 0.37fF


.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create a resistor between the MOSFET drain and VPWR
R VPWR DRAIN 10k

* create pulse
Vin GATE VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10p 2n 0

.control
run
set color0 = white
set color1 = black
plot GATE DRAIN
.endc

.end
