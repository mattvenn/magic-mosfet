magic
tech sky130B
timestamp 1609431046
<< nmos >>
rect 40 0 55 65
<< ndiff >>
rect -5 50 40 65
rect -5 15 0 50
rect 20 15 40 50
rect -5 0 40 15
rect 55 50 100 65
rect 55 15 73 50
rect 93 15 100 50
rect 55 0 100 15
<< ndiffc >>
rect 0 15 20 50
rect 73 15 93 50
<< poly >>
rect 40 65 55 105
rect 40 -10 55 0
rect 15 -25 55 -10
rect 15 -50 20 -25
rect 45 -50 55 -25
rect 15 -58 55 -50
<< polycont >>
rect 20 -50 45 -25
<< locali >>
rect -51 50 26 58
rect -51 49 0 50
rect -51 14 -44 49
rect -25 15 0 49
rect 20 15 26 50
rect -25 14 26 15
rect -51 5 26 14
rect 70 50 147 58
rect 70 15 73 50
rect 93 46 147 50
rect 93 18 115 46
rect 133 18 147 46
rect 93 15 147 18
rect 70 10 147 15
rect 70 5 146 10
rect -25 -23 52 -16
rect -25 -51 -21 -23
rect -3 -25 52 -23
rect -3 -50 20 -25
rect 45 -50 52 -25
rect -3 -51 52 -50
rect -25 -58 52 -51
<< viali >>
rect -44 14 -25 49
rect 115 18 133 46
rect -21 -51 -3 -23
<< metal1 >>
rect -94 49 -12 54
rect -94 14 -44 49
rect -25 14 -12 49
rect -94 11 -12 14
rect 108 46 190 54
rect 108 18 115 46
rect 133 18 190 46
rect 108 11 190 18
rect -80 -23 2 -15
rect -80 -51 -21 -23
rect -3 -51 2 -23
rect -80 -58 2 -51
<< labels >>
rlabel metal1 -90 17 -66 49 1 source
rlabel metal1 -73 -53 -49 -21 1 gate
rlabel metal1 161 15 185 47 1 drain
<< end >>
