* NGSPICE file created from mosfet.ext - technology: sky130A


* Top level circuit mosfet

X0 drain gate source VSUBS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
C0 drain source 0.06fF
C1 gate source 0.20fF
C2 drain VSUBS 0.15fF
C3 source VSUBS 0.15fF
C4 gate VSUBS 0.37fF


