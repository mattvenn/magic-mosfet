magic
tech sky130B
timestamp 1609431327
<< end >>
